module _32bit_2x1MUX(result,A,B,control);
input [31:0] A, B;
input control;
output [31:0] result;

wire [31:0] and1, and2;

and (and1[0], A[0], ~control);
and (and1[1], A[1], ~control);
and (and1[2], A[2], ~control);
and (and1[3], A[3], ~control);
and (and1[4], A[4], ~control);
and (and1[5], A[5], ~control);
and (and1[6], A[6], ~control);
and (and1[7], A[7], ~control);
and (and1[8], A[8], ~control);
and (and1[9], A[9], ~control);
and (and1[10], A[10], ~control);
and (and1[11], A[11], ~control);
and (and1[12], A[12], ~control);
and (and1[13], A[13], ~control);
and (and1[14], A[14], ~control);
and (and1[15], A[15], ~control);
and (and1[16], A[16], ~control);
and (and1[17], A[17], ~control);
and (and1[18], A[18], ~control);
and (and1[19], A[19], ~control);
and (and1[20], A[20], ~control);
and (and1[21], A[21], ~control);
and (and1[22], A[22], ~control);
and (and1[23], A[23], ~control);
and (and1[24], A[24], ~control);
and (and1[25], A[25], ~control);
and (and1[26], A[26], ~control);
and (and1[27], A[27], ~control);
and (and1[28], A[28], ~control);
and (and1[29], A[29], ~control);
and (and1[30], A[30], ~control);
and (and1[31], A[31], ~control);

and (and2[0], B[0], control);
and (and2[1], B[1], control);
and (and2[2], B[2], control);
and (and2[3], B[3], control);
and (and2[4], B[4], control);
and (and2[5], B[5], control);
and (and2[6], B[6], control);
and (and2[7], B[7], control);
and (and2[8], B[8], control);
and (and2[9], B[9], control);
and (and2[10], B[10], control);
and (and2[11], B[11], control);
and (and2[12], B[12], control);
and (and2[13], B[13], control);
and (and2[14], B[14], control);
and (and2[15], B[15], control);
and (and2[16], B[16], control);
and (and2[17], B[17], control);
and (and2[18], B[18], control);
and (and2[19], B[19], control);
and (and2[20], B[20], control);
and (and2[21], B[21], control);
and (and2[22], B[22], control);
and (and2[23], B[23], control);
and (and2[24], B[24], control);
and (and2[25], B[25], control);
and (and2[26], B[26], control);
and (and2[27], B[27], control);
and (and2[28], B[28], control);
and (and2[29], B[29], control);
and (and2[30], B[30], control);
and (and2[31], B[31], control);

or (result[0], and1[0], and2[0]);
or (result[1], and1[1], and2[1]);
or (result[2], and1[2], and2[2]);
or (result[3], and1[3], and2[3]);
or (result[4], and1[4], and2[4]);
or (result[5], and1[5], and2[5]);
or (result[6], and1[6], and2[6]);
or (result[7], and1[7], and2[7]);
or (result[8], and1[8], and2[8]);
or (result[9], and1[9], and2[9]);
or (result[10], and1[10], and2[10]);
or (result[11], and1[11], and2[11]);
or (result[12], and1[12], and2[12]);
or (result[13], and1[13], and2[13]);
or (result[14], and1[14], and2[14]);
or (result[15], and1[15], and2[15]);
or (result[16], and1[16], and2[16]);
or (result[17], and1[17], and2[17]);
or (result[18], and1[18], and2[18]);
or (result[19], and1[19], and2[19]);
or (result[20], and1[20], and2[20]);
or (result[21], and1[21], and2[21]);
or (result[22], and1[22], and2[22]);
or (result[23], and1[23], and2[23]);
or (result[24], and1[24], and2[24]);
or (result[25], and1[25], and2[25]);
or (result[26], and1[26], and2[26]);
or (result[27], and1[27], and2[27]);
or (result[28], and1[28], and2[28]);
or (result[29], and1[29], and2[29]);
or (result[30], and1[30], and2[30]);
or (result[31], and1[31], and2[31]);

endmodule