module spypath_3_1 (N11334, N251, HT_IN1, HT_IN2, Vcc, gnd);
(* keep = 1 *) input HT_IN1, HT_IN2, N251, Vcc, gnd;
(* keep = 1 *) output N11334;
(* keep = 1 *) wire T1, T2, N11313, N11278, N11260, N11321, N11213, N11168, N11115, N11299, N11044, N10988, N10872, N10737, N11328, N10671, N5683, N10672, N6779, N9067, N4471, N1990, N1302, N11242, N3114, N3515, N6783, N9957, N3149, N10989, N10928, N644, N10873, N643, N11314, N6773, N7465, N11114, N6762, N10314, N1833, N8114, N10789, N10509, N10170, N9432, N9066, N10315, N9642, N11214, N9958, N1323, N5171, N7447, N10431, Vcc, gnd;
buf BUFF1_58(N643, N251);
not NOT1_59(N644, N251);
buf BUFF1_162(N1302, N644);
buf BUFF1_169(N1323, N644);
not NOT1_262(N1833, N1302);
and AND2_351(N1990, N644, Vcc);
and AND2_680(N3114, N644, Vcc);
and AND2_691(N3149, N644, Vcc);
nor NOR2_786(N3515, N644, gnd);
nand NAND2_939(N4471, N1833, Vcc);
nand NAND2_1282(N5171, N1302, Vcc);
nand NAND2_1394(N5683, N4471, Vcc);
and AND5_1750(N6762, N5683, Vcc, Vcc, Vcc, Vcc);
and AND4_1758(N6773, N5683, Vcc, Vcc, Vcc);
and AND3_1764(N6779, N5683, Vcc, Vcc);
and AND2_1768(N6783, N5683, Vcc);
buf BUFF1_1959(N7447, N5683);
buf BUFF1_1965(N7465, N5683);
or OR4_2030(N8114, N6779, gnd, gnd, gnd);
not NOT1_2398(N9066, N8114);
nand NAND2_2399(N9067, N8114, Vcc);
nand NAND2_2552(N9432, N9066, Vcc);
nand NAND2_2648(N9642, N9432, Vcc);
not NOT1_2793(N9957, N9642);
nand NAND2_2794(N9958, N9642, Vcc);
nand NAND2_2919(N10170, N9958, Vcc);
not NOT1_2987(N10314, N10170);
nand NAND2_2988(N10315, N10170, Vcc);
nand NAND2_3032(N10431, N10314, Vcc);
nand NAND2_3049(N10509, N10431, Vcc);
not NOT1_3138(N10671, N10509);
nand NAND2_3139(N10672, N10509, Vcc);
nand NAND2_3181(N10737, N10671, Vcc);
nand NAND2_3212(N10789, N10737, Vcc);
not NOT1_3254(N10872, N10789);
nand NAND2_3255(N10873, N10789, Vcc);
nand NAND2_3290(N10928, N10873, Vcc);
not NOT1_3314(N10988, N10928);
nand NAND2_3315(N10989, N10928, Vcc);
nand NAND2_3350(N11044, N10989, Vcc);
not NOT1_3380(N11114, N11044);
nand NAND2_3381(N11115, N11044, Vcc);
nand NAND2_3410(N11168, N11115, Vcc);
not NOT1_3425(N11213, N11168);
nand NAND2_3426(N11214, N11168, Vcc);
nand NAND2_3446(N11242, N11213, Vcc);
nand NAND2_3454(N11260, N11242, Vcc);
and AND2_3466(N11278, N11260, Vcc);
or OR2_3485(N11299, N11278, gnd);
nand NAND2_3491(N11313, N11299, Vcc);
not NOT1_3492(N11314, N11299);

nand HT_TRIGGER(T1, HT_IN1, HT_IN2);
xor HT_PAYLOAD(T2, N11314, T1);

nand NAND2_3497(N11321, T2, Vcc);
nand NAND2_3500(N11328, N11321, Vcc);
not NOT1_3504(N11334, N11328);

endmodule


