module path1(out, in);
input in;
output out;

(* keep = 1 *) wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10,
w11, w12, w13, w14, w15, w16, w17, w18, w19, w20,
w21, w22, w23, w24, w25, w26, w27, w28, w29, w30,
w31, w32, w33, w34, w35, w36, w37, w38, w39, w40,
w41, w42, w43, w44, w45, w46, w47, w48, w49, w50,
w51, w52, w53, w54, w55, w56, w57, w58, w59, w60,
w61, w62, w63, w64, w65, w66, w67, w68, w69, w70,
w71, w72, w73, w74, w75, w76, w77, w78, w79, w80,
w81, w82, w83, w84, w85, w86, w87, w88, w89, w90,
w91, w92, w93, w94, w95, w96, w97, w98, w99, w100,
w101, w102, w103, w104, w105, w106, w107, w108, w109, w110,
w111, w112, w113, w114, w115, w116, w117, w118, w119, w120,
w121, w122, w123, w124, w125, w126, w127, w128, w129, w130,
w131, w132, w133, w134, w135, w136, w137, w138, w139, w140,
w141, w142, w143, w144, w145, w146, w147, w148, w149, w150,
w151, w152, w153, w154, w155, w156, w157, w158, w159, w160,
w161, w162, w163, w164, w165, w166, w167, w168, w169, w170,
w171, w172, w173, w174, w175, w176, w177, w178, w179, w180,
w181, w182, w183, w184, w185, w186, w187, w188, w189, w190,
w191, w192, w193, w194, w195, w196, w197, w198, w199, w200,
w201, w202, w203, w204, w205, w206, w207, w208, w209, w210,
w211, w212, w213, w214, w215, w216, w217, w218, w219, w220,
w221, w222, w223, w224, w225, w226, w227, w228, w229, w230,
w231, w232, w233, w234, w235, w236, w237, w238, w239, w240,
w241, w242, w243, w244, w245, w246, w247, w248, w249, w250,
w251, w252, w253, w254, w255, w256, w257, w258, w259, w260,
w261, w262, w263, w264, w265, w266, w267, w268, w269, w270,
w271, w272, w273, w274, w275, w276, w277, w278, w279, w280,
w281, w282, w283, w284, w285, w286, w287, w288, w289, w290,
w291, w292, w293, w294, w295, w296, w297, w298, w299, w300,
w301, w302, w303, w304, w305, w306, w307, w308, w309, w310,
w311, w312, w313, w314, w315, w316, w317, w318, w319, w320,
w321, w322, w323, w324, w325, w326, w327, w328, w329, w330,
w331, w332, w333, w334, w335, w336, w337, w338, w339, w340,
w341, w342, w343, w344, w345, w346, w347, w348, w349, w350,
w351, w352, w353, w354, w355, w356, w357, w358, w359, w360,
w361, w362, w363, w364, w365, w366, w367, w368, w369, w370,
w371, w372, w373, w374, w375, w376, w377, w378, w379, w380,
w381, w382, w383, w384, w385, w386, w387, w388, w389, w390,
w391, w392, w393, w394, w395, w396, w397, w398, w399, w400,
w401, w402, w403, w404, w405, w406, w407, w408, w409, w410,
w411, w412, w413, w414, w415, w416, w417, w418, w419, w420,
w421, w422, w423, w424, w425, w426, w427, w428, w429, w430,
w431, w432, w433, w434, w435, w436, w437, w438, w439, w440,
w441, w442, w443, w444, w445, w446, w447, w448, w449, w450,
w451, w452, w453, w454, w455, w456, w457, w458, w459, w460,
w461, w462, w463, w464, w465, w466, w467, w468, w469, w470,
w471, w472, w473, w474, w475, w476, w477, w478, w479, w480,
w481, w482, w483, w484, w485, w486, w487, w488, w489, w490,
w491, w492, w493, w494, w495, w496, w497, w498, w499, w500,
w501, w502, w503, w504, w505, w506, w507, w508, w509, w510,
w511, w512, w513, w514, w515, w516, w517, w518, w519, w520,
w521, w522, w523, w524, w525, w526, w527, w528, w529, w530,
w531, w532, w533, w534, w535, w536, w537, w538, w539, w540,
w541, w542, w543, w544, w545, w546, w547, w548, w549, w550,
w551, w552, w553, w554, w555, w556, w557, w558, w559, w560,
w561, w562, w563, w564, w565, w566, w567, w568, w569, w570,
w571, w572, w573, w574, w575, w576, w577, w578, w579, w580,
w581, w582, w583, w584, w585, w586, w587, w588, w589, w590,
w591, w592, w593, w594, w595, w596, w597, w598, w599, w600,
w601, w602, w603, w604, w605, w606, w607, w608, w609, w610,
w611, w612, w613, w614, w615, w616, w617, w618, w619, w620,
w621, w622, w623, w624, w625, w626, w627, w628, w629, w630,
w631, w632, w633, w634, w635, w636, w637, w638, w639, w640,
w641, w642, w643, w644, w645, w646, w647, w648, w649, w650,
w651, w652, w653, w654, w655, w656, w657, w658, w659, w660,
w661, w662, w663, w664, w665, w666, w667, w668, w669, w670,
w671, w672, w673, w674, w675, w676, w677, w678, w679, w680,
w681, w682, w683, w684, w685, w686, w687, w688, w689, w690,
w691, w692, w693, w694, w695, w696, w697, w698, w699, w700,
w701, w702, w703, w704, w705, w706, w707, w708, w709, w710,
w711, w712, w713, w714, w715, w716, w717, w718, w719, w720,
w721, w722, w723, w724, w725, w726, w727, w728, w729, w730,
w731, w732, w733, w734, w735, w736, w737, w738, w739, w740,
w741, w742, w743, w744, w745, w746, w747, w748, w749, w750,
w751, w752, w753, w754, w755, w756, w757, w758, w759, w760,
w761, w762, w763, w764, w765, w766, w767, w768, w769, w770,
w771, w772, w773, w774, w775, w776, w777, w778, w779, w780,
w781, w782, w783, w784, w785, w786, w787, w788, w789, w790,
w791, w792, w793, w794, w795, w796, w797, w798, w799, w800,
w801, w802, w803, w804, w805, w806, w807, w808, w809, w810,
w811, w812, w813, w814, w815, w816, w817, w818, w819, w820,
w821, w822, w823, w824, w825, w826, w827, w828, w829, w830,
w831, w832, w833, w834, w835, w836, w837, w838, w839, w840,
w841, w842, w843, w844, w845, w846, w847, w848, w849, w850,
w851, w852, w853, w854, w855, w856, w857, w858, w859, w860,
w861, w862, w863, w864, w865, w866, w867, w868, w869, w870,
w871, w872, w873, w874, w875, w876, w877, w878, w879, w880,
w881, w882, w883, w884, w885, w886, w887, w888, w889, w890,
w891, w892, w893, w894, w895, w896, w897, w898, w899, w900,
w901, w902, w903, w904, w905, w906, w907, w908, w909, w910,
w911, w912, w913, w914, w915, w916, w917, w918, w919, w920,
w921, w922, w923, w924, w925, w926, w927, w928, w929, w930,
w931, w932, w933, w934, w935, w936, w937, w938, w939, w940,
w941, w942, w943, w944, w945, w946, w947, w948, w949, w950,
w951, w952, w953, w954, w955, w956, w957, w958, w959, w960,
w961, w962, w963, w964, w965, w966, w967, w968, w969, w970,
w971, w972, w973, w974, w975, w976, w977, w978, w979, w980,
w981, w982, w983, w984, w985, w986, w987, w988, w989, w990,
w991, w992, w993, w994, w995, w996, w997, w998;

not n0(w0, in);
not n1(w1, w0);
not n2(w2, w1);
not n3(w3, w2);
not n4(w4, w3);
not n5(w5, w4);
not n6(w6, w5);
not n7(w7, w6);
not n8(w8, w7);
not n9(w9, w8);
not n10(w10, w9);
not n11(w11, w10);
not n12(w12, w11);
not n13(w13, w12);
not n14(w14, w13);
not n15(w15, w14);
not n16(w16, w15);
not n17(w17, w16);
not n18(w18, w17);
not n19(w19, w18);
not n20(w20, w19);
not n21(w21, w20);
not n22(w22, w21);
not n23(w23, w22);
not n24(w24, w23);
not n25(w25, w24);
not n26(w26, w25);
not n27(w27, w26);
not n28(w28, w27);
not n29(w29, w28);
not n30(w30, w29);
not n31(w31, w30);
not n32(w32, w31);
not n33(w33, w32);
not n34(w34, w33);
not n35(w35, w34);
not n36(w36, w35);
not n37(w37, w36);
not n38(w38, w37);
not n39(w39, w38);
not n40(w40, w39);
not n41(w41, w40);
not n42(w42, w41);
not n43(w43, w42);
not n44(w44, w43);
not n45(w45, w44);
not n46(w46, w45);
not n47(w47, w46);
not n48(w48, w47);
not n49(w49, w48);
not n50(w50, w49);
not n51(w51, w50);
not n52(w52, w51);
not n53(w53, w52);
not n54(w54, w53);
not n55(w55, w54);
not n56(w56, w55);
not n57(w57, w56);
not n58(w58, w57);
not n59(w59, w58);
not n60(w60, w59);
not n61(w61, w60);
not n62(w62, w61);
not n63(w63, w62);
not n64(w64, w63);
not n65(w65, w64);
not n66(w66, w65);
not n67(w67, w66);
not n68(w68, w67);
not n69(w69, w68);
not n70(w70, w69);
not n71(w71, w70);
not n72(w72, w71);
not n73(w73, w72);
not n74(w74, w73);
not n75(w75, w74);
not n76(w76, w75);
not n77(w77, w76);
not n78(w78, w77);
not n79(w79, w78);
not n80(w80, w79);
not n81(w81, w80);
not n82(w82, w81);
not n83(w83, w82);
not n84(w84, w83);
not n85(w85, w84);
not n86(w86, w85);
not n87(w87, w86);
not n88(w88, w87);
not n89(w89, w88);
not n90(w90, w89);
not n91(w91, w90);
not n92(w92, w91);
not n93(w93, w92);
not n94(w94, w93);
not n95(w95, w94);
not n96(w96, w95);
not n97(w97, w96);
not n98(w98, w97);
not n99(w99, w98);
not n100(w100, w99);
not n101(w101, w100);
not n102(w102, w101);
not n103(w103, w102);
not n104(w104, w103);
not n105(w105, w104);
not n106(w106, w105);
not n107(w107, w106);
not n108(w108, w107);
not n109(w109, w108);
not n110(w110, w109);
not n111(w111, w110);
not n112(w112, w111);
not n113(w113, w112);
not n114(w114, w113);
not n115(w115, w114);
not n116(w116, w115);
not n117(w117, w116);
not n118(w118, w117);
not n119(w119, w118);
not n120(w120, w119);
not n121(w121, w120);
not n122(w122, w121);
not n123(w123, w122);
not n124(w124, w123);
not n125(w125, w124);
not n126(w126, w125);
not n127(w127, w126);
not n128(w128, w127);
not n129(w129, w128);
not n130(w130, w129);
not n131(w131, w130);
not n132(w132, w131);
not n133(w133, w132);
not n134(w134, w133);
not n135(w135, w134);
not n136(w136, w135);
not n137(w137, w136);
not n138(w138, w137);
not n139(w139, w138);
not n140(w140, w139);
not n141(w141, w140);
not n142(w142, w141);
not n143(w143, w142);
not n144(w144, w143);
not n145(w145, w144);
not n146(w146, w145);
not n147(w147, w146);
not n148(w148, w147);
not n149(w149, w148);
not n150(w150, w149);
not n151(w151, w150);
not n152(w152, w151);
not n153(w153, w152);
not n154(w154, w153);
not n155(w155, w154);
not n156(w156, w155);
not n157(w157, w156);
not n158(w158, w157);
not n159(w159, w158);
not n160(w160, w159);
not n161(w161, w160);
not n162(w162, w161);
not n163(w163, w162);
not n164(w164, w163);
not n165(w165, w164);
not n166(w166, w165);
not n167(w167, w166);
not n168(w168, w167);
not n169(w169, w168);
not n170(w170, w169);
not n171(w171, w170);
not n172(w172, w171);
not n173(w173, w172);
not n174(w174, w173);
not n175(w175, w174);
not n176(w176, w175);
not n177(w177, w176);
not n178(w178, w177);
not n179(w179, w178);
not n180(w180, w179);
not n181(w181, w180);
not n182(w182, w181);
not n183(w183, w182);
not n184(w184, w183);
not n185(w185, w184);
not n186(w186, w185);
not n187(w187, w186);
not n188(w188, w187);
not n189(w189, w188);
not n190(w190, w189);
not n191(w191, w190);
not n192(w192, w191);
not n193(w193, w192);
not n194(w194, w193);
not n195(w195, w194);
not n196(w196, w195);
not n197(w197, w196);
not n198(w198, w197);
not n199(w199, w198);
not n200(w200, w199);
not n201(w201, w200);
not n202(w202, w201);
not n203(w203, w202);
not n204(w204, w203);
not n205(w205, w204);
not n206(w206, w205);
not n207(w207, w206);
not n208(w208, w207);
not n209(w209, w208);
not n210(w210, w209);
not n211(w211, w210);
not n212(w212, w211);
not n213(w213, w212);
not n214(w214, w213);
not n215(w215, w214);
not n216(w216, w215);
not n217(w217, w216);
not n218(w218, w217);
not n219(w219, w218);
not n220(w220, w219);
not n221(w221, w220);
not n222(w222, w221);
not n223(w223, w222);
not n224(w224, w223);
not n225(w225, w224);
not n226(w226, w225);
not n227(w227, w226);
not n228(w228, w227);
not n229(w229, w228);
not n230(w230, w229);
not n231(w231, w230);
not n232(w232, w231);
not n233(w233, w232);
not n234(w234, w233);
not n235(w235, w234);
not n236(w236, w235);
not n237(w237, w236);
not n238(w238, w237);
not n239(w239, w238);
not n240(w240, w239);
not n241(w241, w240);
not n242(w242, w241);
not n243(w243, w242);
not n244(w244, w243);
not n245(w245, w244);
not n246(w246, w245);
not n247(w247, w246);
not n248(w248, w247);
not n249(w249, w248);
not n250(w250, w249);
not n251(w251, w250);
not n252(w252, w251);
not n253(w253, w252);
not n254(w254, w253);
not n255(w255, w254);
not n256(w256, w255);
not n257(w257, w256);
not n258(w258, w257);
not n259(w259, w258);
not n260(w260, w259);
not n261(w261, w260);
not n262(w262, w261);
not n263(w263, w262);
not n264(w264, w263);
not n265(w265, w264);
not n266(w266, w265);
not n267(w267, w266);
not n268(w268, w267);
not n269(w269, w268);
not n270(w270, w269);
not n271(w271, w270);
not n272(w272, w271);
not n273(w273, w272);
not n274(w274, w273);
not n275(w275, w274);
not n276(w276, w275);
not n277(w277, w276);
not n278(w278, w277);
not n279(w279, w278);
not n280(w280, w279);
not n281(w281, w280);
not n282(w282, w281);
not n283(w283, w282);
not n284(w284, w283);
not n285(w285, w284);
not n286(w286, w285);
not n287(w287, w286);
not n288(w288, w287);
not n289(w289, w288);
not n290(w290, w289);
not n291(w291, w290);
not n292(w292, w291);
not n293(w293, w292);
not n294(w294, w293);
not n295(w295, w294);
not n296(w296, w295);
not n297(w297, w296);
not n298(w298, w297);
not n299(w299, w298);
not n300(w300, w299);
not n301(w301, w300);
not n302(w302, w301);
not n303(w303, w302);
not n304(w304, w303);
not n305(w305, w304);
not n306(w306, w305);
not n307(w307, w306);
not n308(w308, w307);
not n309(w309, w308);
not n310(w310, w309);
not n311(w311, w310);
not n312(w312, w311);
not n313(w313, w312);
not n314(w314, w313);
not n315(w315, w314);
not n316(w316, w315);
not n317(w317, w316);
not n318(w318, w317);
not n319(w319, w318);
not n320(w320, w319);
not n321(w321, w320);
not n322(w322, w321);
not n323(w323, w322);
not n324(w324, w323);
not n325(w325, w324);
not n326(w326, w325);
not n327(w327, w326);
not n328(w328, w327);
not n329(w329, w328);
not n330(w330, w329);
not n331(w331, w330);
not n332(w332, w331);
not n333(w333, w332);
not n334(w334, w333);
not n335(w335, w334);
not n336(w336, w335);
not n337(w337, w336);
not n338(w338, w337);
not n339(w339, w338);
not n340(w340, w339);
not n341(w341, w340);
not n342(w342, w341);
not n343(w343, w342);
not n344(w344, w343);
not n345(w345, w344);
not n346(w346, w345);
not n347(w347, w346);
not n348(w348, w347);
not n349(w349, w348);
not n350(w350, w349);
not n351(w351, w350);
not n352(w352, w351);
not n353(w353, w352);
not n354(w354, w353);
not n355(w355, w354);
not n356(w356, w355);
not n357(w357, w356);
not n358(w358, w357);
not n359(w359, w358);
not n360(w360, w359);
not n361(w361, w360);
not n362(w362, w361);
not n363(w363, w362);
not n364(w364, w363);
not n365(w365, w364);
not n366(w366, w365);
not n367(w367, w366);
not n368(w368, w367);
not n369(w369, w368);
not n370(w370, w369);
not n371(w371, w370);
not n372(w372, w371);
not n373(w373, w372);
not n374(w374, w373);
not n375(w375, w374);
not n376(w376, w375);
not n377(w377, w376);
not n378(w378, w377);
not n379(w379, w378);
not n380(w380, w379);
not n381(w381, w380);
not n382(w382, w381);
not n383(w383, w382);
not n384(w384, w383);
not n385(w385, w384);
not n386(w386, w385);
not n387(w387, w386);
not n388(w388, w387);
not n389(w389, w388);
not n390(w390, w389);
not n391(w391, w390);
not n392(w392, w391);
not n393(w393, w392);
not n394(w394, w393);
not n395(w395, w394);
not n396(w396, w395);
not n397(w397, w396);
not n398(w398, w397);
not n399(w399, w398);
not n400(w400, w399);
not n401(w401, w400);
not n402(w402, w401);
not n403(w403, w402);
not n404(w404, w403);
not n405(w405, w404);
not n406(w406, w405);
not n407(w407, w406);
not n408(w408, w407);
not n409(w409, w408);
not n410(w410, w409);
not n411(w411, w410);
not n412(w412, w411);
not n413(w413, w412);
not n414(w414, w413);
not n415(w415, w414);
not n416(w416, w415);
not n417(w417, w416);
not n418(w418, w417);
not n419(w419, w418);
not n420(w420, w419);
not n421(w421, w420);
not n422(w422, w421);
not n423(w423, w422);
not n424(w424, w423);
not n425(w425, w424);
not n426(w426, w425);
not n427(w427, w426);
not n428(w428, w427);
not n429(w429, w428);
not n430(w430, w429);
not n431(w431, w430);
not n432(w432, w431);
not n433(w433, w432);
not n434(w434, w433);
not n435(w435, w434);
not n436(w436, w435);
not n437(w437, w436);
not n438(w438, w437);
not n439(w439, w438);
not n440(w440, w439);
not n441(w441, w440);
not n442(w442, w441);
not n443(w443, w442);
not n444(w444, w443);
not n445(w445, w444);
not n446(w446, w445);
not n447(w447, w446);
not n448(w448, w447);
not n449(w449, w448);
not n450(w450, w449);
not n451(w451, w450);
not n452(w452, w451);
not n453(w453, w452);
not n454(w454, w453);
not n455(w455, w454);
not n456(w456, w455);
not n457(w457, w456);
not n458(w458, w457);
not n459(w459, w458);
not n460(w460, w459);
not n461(w461, w460);
not n462(w462, w461);
not n463(w463, w462);
not n464(w464, w463);
not n465(w465, w464);
not n466(w466, w465);
not n467(w467, w466);
not n468(w468, w467);
not n469(w469, w468);
not n470(w470, w469);
not n471(w471, w470);
not n472(w472, w471);
not n473(w473, w472);
not n474(w474, w473);
not n475(w475, w474);
not n476(w476, w475);
not n477(w477, w476);
not n478(w478, w477);
not n479(w479, w478);
not n480(w480, w479);
not n481(w481, w480);
not n482(w482, w481);
not n483(w483, w482);
not n484(w484, w483);
not n485(w485, w484);
not n486(w486, w485);
not n487(w487, w486);
not n488(w488, w487);
not n489(w489, w488);
not n490(w490, w489);
not n491(w491, w490);
not n492(w492, w491);
not n493(w493, w492);
not n494(w494, w493);
not n495(w495, w494);
not n496(w496, w495);
not n497(w497, w496);
not n498(w498, w497);
not n499(w499, w498);
not n500(w500, w499);
not n501(w501, w500);
not n502(w502, w501);
not n503(w503, w502);
not n504(w504, w503);
not n505(w505, w504);
not n506(w506, w505);
not n507(w507, w506);
not n508(w508, w507);
not n509(w509, w508);
not n510(w510, w509);
not n511(w511, w510);
not n512(w512, w511);
not n513(w513, w512);
not n514(w514, w513);
not n515(w515, w514);
not n516(w516, w515);
not n517(w517, w516);
not n518(w518, w517);
not n519(w519, w518);
not n520(w520, w519);
not n521(w521, w520);
not n522(w522, w521);
not n523(w523, w522);
not n524(w524, w523);
not n525(w525, w524);
not n526(w526, w525);
not n527(w527, w526);
not n528(w528, w527);
not n529(w529, w528);
not n530(w530, w529);
not n531(w531, w530);
not n532(w532, w531);
not n533(w533, w532);
not n534(w534, w533);
not n535(w535, w534);
not n536(w536, w535);
not n537(w537, w536);
not n538(w538, w537);
not n539(w539, w538);
not n540(w540, w539);
not n541(w541, w540);
not n542(w542, w541);
not n543(w543, w542);
not n544(w544, w543);
not n545(w545, w544);
not n546(w546, w545);
not n547(w547, w546);
not n548(w548, w547);
not n549(w549, w548);
not n550(w550, w549);
not n551(w551, w550);
not n552(w552, w551);
not n553(w553, w552);
not n554(w554, w553);
not n555(w555, w554);
not n556(w556, w555);
not n557(w557, w556);
not n558(w558, w557);
not n559(w559, w558);
not n560(w560, w559);
not n561(w561, w560);
not n562(w562, w561);
not n563(w563, w562);
not n564(w564, w563);
not n565(w565, w564);
not n566(w566, w565);
not n567(w567, w566);
not n568(w568, w567);
not n569(w569, w568);
not n570(w570, w569);
not n571(w571, w570);
not n572(w572, w571);
not n573(w573, w572);
not n574(w574, w573);
not n575(w575, w574);
not n576(w576, w575);
not n577(w577, w576);
not n578(w578, w577);
not n579(w579, w578);
not n580(w580, w579);
not n581(w581, w580);
not n582(w582, w581);
not n583(w583, w582);
not n584(w584, w583);
not n585(w585, w584);
not n586(w586, w585);
not n587(w587, w586);
not n588(w588, w587);
not n589(w589, w588);
not n590(w590, w589);
not n591(w591, w590);
not n592(w592, w591);
not n593(w593, w592);
not n594(w594, w593);
not n595(w595, w594);
not n596(w596, w595);
not n597(w597, w596);
not n598(w598, w597);
not n599(w599, w598);
not n600(w600, w599);
not n601(w601, w600);
not n602(w602, w601);
not n603(w603, w602);
not n604(w604, w603);
not n605(w605, w604);
not n606(w606, w605);
not n607(w607, w606);
not n608(w608, w607);
not n609(w609, w608);
not n610(w610, w609);
not n611(w611, w610);
not n612(w612, w611);
not n613(w613, w612);
not n614(w614, w613);
not n615(w615, w614);
not n616(w616, w615);
not n617(w617, w616);
not n618(w618, w617);
not n619(w619, w618);
not n620(w620, w619);
not n621(w621, w620);
not n622(w622, w621);
not n623(w623, w622);
not n624(w624, w623);
not n625(w625, w624);
not n626(w626, w625);
not n627(w627, w626);
not n628(w628, w627);
not n629(w629, w628);
not n630(w630, w629);
not n631(w631, w630);
not n632(w632, w631);
not n633(w633, w632);
not n634(w634, w633);
not n635(w635, w634);
not n636(w636, w635);
not n637(w637, w636);
not n638(w638, w637);
not n639(w639, w638);
not n640(w640, w639);
not n641(w641, w640);
not n642(w642, w641);
not n643(w643, w642);
not n644(w644, w643);
not n645(w645, w644);
not n646(w646, w645);
not n647(w647, w646);
not n648(w648, w647);
not n649(w649, w648);
not n650(w650, w649);
not n651(w651, w650);
not n652(w652, w651);
not n653(w653, w652);
not n654(w654, w653);
not n655(w655, w654);
not n656(w656, w655);
not n657(w657, w656);
not n658(w658, w657);
not n659(w659, w658);
not n660(w660, w659);
not n661(w661, w660);
not n662(w662, w661);
not n663(w663, w662);
not n664(w664, w663);
not n665(w665, w664);
not n666(w666, w665);
not n667(w667, w666);
not n668(w668, w667);
not n669(w669, w668);
not n670(w670, w669);
not n671(w671, w670);
not n672(w672, w671);
not n673(w673, w672);
not n674(w674, w673);
not n675(w675, w674);
not n676(w676, w675);
not n677(w677, w676);
not n678(w678, w677);
not n679(w679, w678);
not n680(w680, w679);
not n681(w681, w680);
not n682(w682, w681);
not n683(w683, w682);
not n684(w684, w683);
not n685(w685, w684);
not n686(w686, w685);
not n687(w687, w686);
not n688(w688, w687);
not n689(w689, w688);
not n690(w690, w689);
not n691(w691, w690);
not n692(w692, w691);
not n693(w693, w692);
not n694(w694, w693);
not n695(w695, w694);
not n696(w696, w695);
not n697(w697, w696);
not n698(w698, w697);
not n699(w699, w698);
not n700(w700, w699);
not n701(w701, w700);
not n702(w702, w701);
not n703(w703, w702);
not n704(w704, w703);
not n705(w705, w704);
not n706(w706, w705);
not n707(w707, w706);
not n708(w708, w707);
not n709(w709, w708);
not n710(w710, w709);
not n711(w711, w710);
not n712(w712, w711);
not n713(w713, w712);
not n714(w714, w713);
not n715(w715, w714);
not n716(w716, w715);
not n717(w717, w716);
not n718(w718, w717);
not n719(w719, w718);
not n720(w720, w719);
not n721(w721, w720);
not n722(w722, w721);
not n723(w723, w722);
not n724(w724, w723);
not n725(w725, w724);
not n726(w726, w725);
not n727(w727, w726);
not n728(w728, w727);
not n729(w729, w728);
not n730(w730, w729);
not n731(w731, w730);
not n732(w732, w731);
not n733(w733, w732);
not n734(w734, w733);
not n735(w735, w734);
not n736(w736, w735);
not n737(w737, w736);
not n738(w738, w737);
not n739(w739, w738);
not n740(w740, w739);
not n741(w741, w740);
not n742(w742, w741);
not n743(w743, w742);
not n744(w744, w743);
not n745(w745, w744);
not n746(w746, w745);
not n747(w747, w746);
not n748(w748, w747);
not n749(w749, w748);
not n750(w750, w749);
not n751(w751, w750);
not n752(w752, w751);
not n753(w753, w752);
not n754(w754, w753);
not n755(w755, w754);
not n756(w756, w755);
not n757(w757, w756);
not n758(w758, w757);
not n759(w759, w758);
not n760(w760, w759);
not n761(w761, w760);
not n762(w762, w761);
not n763(w763, w762);
not n764(w764, w763);
not n765(w765, w764);
not n766(w766, w765);
not n767(w767, w766);
not n768(w768, w767);
not n769(w769, w768);
not n770(w770, w769);
not n771(w771, w770);
not n772(w772, w771);
not n773(w773, w772);
not n774(w774, w773);
not n775(w775, w774);
not n776(w776, w775);
not n777(w777, w776);
not n778(w778, w777);
not n779(w779, w778);
not n780(w780, w779);
not n781(w781, w780);
not n782(w782, w781);
not n783(w783, w782);
not n784(w784, w783);
not n785(w785, w784);
not n786(w786, w785);
not n787(w787, w786);
not n788(w788, w787);
not n789(w789, w788);
not n790(w790, w789);
not n791(w791, w790);
not n792(w792, w791);
not n793(w793, w792);
not n794(w794, w793);
not n795(w795, w794);
not n796(w796, w795);
not n797(w797, w796);
not n798(w798, w797);
not n799(w799, w798);
not n800(w800, w799);
not n801(w801, w800);
not n802(w802, w801);
not n803(w803, w802);
not n804(w804, w803);
not n805(w805, w804);
not n806(w806, w805);
not n807(w807, w806);
not n808(w808, w807);
not n809(w809, w808);
not n810(w810, w809);
not n811(w811, w810);
not n812(w812, w811);
not n813(w813, w812);
not n814(w814, w813);
not n815(w815, w814);
not n816(w816, w815);
not n817(w817, w816);
not n818(w818, w817);
not n819(w819, w818);
not n820(w820, w819);
not n821(w821, w820);
not n822(w822, w821);
not n823(w823, w822);
not n824(w824, w823);
not n825(w825, w824);
not n826(w826, w825);
not n827(w827, w826);
not n828(w828, w827);
not n829(w829, w828);
not n830(w830, w829);
not n831(w831, w830);
not n832(w832, w831);
not n833(w833, w832);
not n834(w834, w833);
not n835(w835, w834);
not n836(w836, w835);
not n837(w837, w836);
not n838(w838, w837);
not n839(w839, w838);
not n840(w840, w839);
not n841(w841, w840);
not n842(w842, w841);
not n843(w843, w842);
not n844(w844, w843);
not n845(w845, w844);
not n846(w846, w845);
not n847(w847, w846);
not n848(w848, w847);
not n849(w849, w848);
not n850(w850, w849);
not n851(w851, w850);
not n852(w852, w851);
not n853(w853, w852);
not n854(w854, w853);
not n855(w855, w854);
not n856(w856, w855);
not n857(w857, w856);
not n858(w858, w857);
not n859(w859, w858);
not n860(w860, w859);
not n861(w861, w860);
not n862(w862, w861);
not n863(w863, w862);
not n864(w864, w863);
not n865(w865, w864);
not n866(w866, w865);
not n867(w867, w866);
not n868(w868, w867);
not n869(w869, w868);
not n870(w870, w869);
not n871(w871, w870);
not n872(w872, w871);
not n873(w873, w872);
not n874(w874, w873);
not n875(w875, w874);
not n876(w876, w875);
not n877(w877, w876);
not n878(w878, w877);
not n879(w879, w878);
not n880(w880, w879);
not n881(w881, w880);
not n882(w882, w881);
not n883(w883, w882);
not n884(w884, w883);
not n885(w885, w884);
not n886(w886, w885);
not n887(w887, w886);
not n888(w888, w887);
not n889(w889, w888);
not n890(w890, w889);
not n891(w891, w890);
not n892(w892, w891);
not n893(w893, w892);
not n894(w894, w893);
not n895(w895, w894);
not n896(w896, w895);
not n897(w897, w896);
not n898(w898, w897);
not n899(w899, w898);
not n900(w900, w899);
not n901(w901, w900);
not n902(w902, w901);
not n903(w903, w902);
not n904(w904, w903);
not n905(w905, w904);
not n906(w906, w905);
not n907(w907, w906);
not n908(w908, w907);
not n909(w909, w908);
not n910(w910, w909);
not n911(w911, w910);
not n912(w912, w911);
not n913(w913, w912);
not n914(w914, w913);
not n915(w915, w914);
not n916(w916, w915);
not n917(w917, w916);
not n918(w918, w917);
not n919(w919, w918);
not n920(w920, w919);
not n921(w921, w920);
not n922(w922, w921);
not n923(w923, w922);
not n924(w924, w923);
not n925(w925, w924);
not n926(w926, w925);
not n927(w927, w926);
not n928(w928, w927);
not n929(w929, w928);
not n930(w930, w929);
not n931(w931, w930);
not n932(w932, w931);
not n933(w933, w932);
not n934(w934, w933);
not n935(w935, w934);
not n936(w936, w935);
not n937(w937, w936);
not n938(w938, w937);
not n939(w939, w938);
not n940(w940, w939);
not n941(w941, w940);
not n942(w942, w941);
not n943(w943, w942);
not n944(w944, w943);
not n945(w945, w944);
not n946(w946, w945);
not n947(w947, w946);
not n948(w948, w947);
not n949(w949, w948);
not n950(w950, w949);
not n951(w951, w950);
not n952(w952, w951);
not n953(w953, w952);
not n954(w954, w953);
not n955(w955, w954);
not n956(w956, w955);
not n957(w957, w956);
not n958(w958, w957);
not n959(w959, w958);
not n960(w960, w959);
not n961(w961, w960);
not n962(w962, w961);
not n963(w963, w962);
not n964(w964, w963);
not n965(w965, w964);
not n966(w966, w965);
not n967(w967, w966);
not n968(w968, w967);
not n969(w969, w968);
not n970(w970, w969);
not n971(w971, w970);
not n972(w972, w971);
not n973(w973, w972);
not n974(w974, w973);
not n975(w975, w974);
not n976(w976, w975);
not n977(w977, w976);
not n978(w978, w977);
not n979(w979, w978);
not n980(w980, w979);
not n981(w981, w980);
not n982(w982, w981);
not n983(w983, w982);
not n984(w984, w983);
not n985(w985, w984);
not n986(w986, w985);
not n987(w987, w986);
not n988(w988, w987);
not n989(w989, w988);
not n990(w990, w989);
not n991(w991, w990);
not n992(w992, w991);
not n993(w993, w992);
not n994(w994, w993);
not n995(w995, w994);
not n996(w996, w995);
not n997(w997, w996);
not n998(w998, w997);
not n999(out, w998);
endmodule
